class Transaction;
	rand bit[2:0]in1;
	rand bit[2:0]in2;
	bit clk;
	bit[3:0]out;	
endclass